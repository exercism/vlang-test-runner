module main

fn is_leap_year123BahB214